// tb_projection_inst.v

// Generated using ACDS version 21.1 850

`timescale 1 ps / 1 ps
module tb_projection_inst (
		input  wire         start,                  //             call.valid
		output wire         busy,                   //                 .stall
		input  wire         clock,                  //            clock.clk
		input  wire         resetn,                 //            reset.reset_n
		output wire         done,                   //           return.valid
		input  wire         stall,                  //                 .stall
		input  wire [351:0] stream_in_tuple_data,   //  stream_in_tuple.data
		output wire         stream_in_tuple_ready,  //                 .ready
		input  wire         stream_in_tuple_valid,  //                 .valid
		output wire [351:0] stream_out_tuple_data,  // stream_out_tuple.data
		input  wire         stream_out_tuple_ready, //                 .ready
		output wire         stream_out_tuple_valid  //                 .valid
	);

	projection_internal projection_internal_inst (
		.clock                  (clock),                  //            clock.clk
		.resetn                 (resetn),                 //            reset.reset_n
		.stream_in_tuple_data   (stream_in_tuple_data),   //  stream_in_tuple.data
		.stream_in_tuple_ready  (stream_in_tuple_ready),  //                 .ready
		.stream_in_tuple_valid  (stream_in_tuple_valid),  //                 .valid
		.stream_out_tuple_data  (stream_out_tuple_data),  // stream_out_tuple.data
		.stream_out_tuple_ready (stream_out_tuple_ready), //                 .ready
		.stream_out_tuple_valid (stream_out_tuple_valid), //                 .valid
		.start                  (start),                  //             call.valid
		.busy                   (busy),                   //                 .stall
		.done                   (done),                   //           return.valid
		.stall                  (stall)                   //                 .stall
	);

endmodule
