// tb.v

// Generated using ACDS version 21.1 850

`timescale 1 ps / 1 ps
module tb (
	);

	wire          streamer_inst_s_out_valid;                                                            // streamer_inst:s_out_valid -> stream_sink_dpi_bfm_streamer_s_out_inst:sink_valid
	wire  [351:0] streamer_inst_s_out_data;                                                             // streamer_inst:s_out_data -> stream_sink_dpi_bfm_streamer_s_out_inst:sink_data
	wire          streamer_inst_s_out_ready;                                                            // stream_sink_dpi_bfm_streamer_s_out_inst:sink_ready -> streamer_inst:s_out_ready
	wire          stream_source_dpi_bfm_streamer_s_in_inst_source_valid;                                // stream_source_dpi_bfm_streamer_s_in_inst:source_valid -> streamer_inst:s_in_valid
	wire  [351:0] stream_source_dpi_bfm_streamer_s_in_inst_source_data;                                 // stream_source_dpi_bfm_streamer_s_in_inst:source_data -> streamer_inst:s_in_data
	wire          stream_source_dpi_bfm_streamer_s_in_inst_source_ready;                                // streamer_inst:s_in_ready -> stream_source_dpi_bfm_streamer_s_in_inst:source_ready
	wire          clock_reset_inst_clock_clk;                                                           // clock_reset_inst:clock -> [component_dpi_controller_streamer_inst:clock, irq_mapper:clk, main_dpi_controller_inst:clock, stream_sink_dpi_bfm_streamer_s_out_inst:clock, stream_source_dpi_bfm_streamer_s_in_inst:clock, streamer_inst:clock]
	wire          clock_reset_inst_clock2x_clk;                                                         // clock_reset_inst:clock2x -> [component_dpi_controller_streamer_inst:clock2x, main_dpi_controller_inst:clock2x, stream_sink_dpi_bfm_streamer_s_out_inst:clock2x, stream_source_dpi_bfm_streamer_s_in_inst:clock2x]
	wire          component_dpi_controller_streamer_inst_component_call_valid;                          // component_dpi_controller_streamer_inst:start -> streamer_inst:start
	wire          streamer_inst_call_stall;                                                             // streamer_inst:busy -> component_dpi_controller_streamer_inst:busy
	wire          component_dpi_controller_streamer_inst_component_done_conduit;                        // component_dpi_controller_streamer_inst:component_done -> concatenate_component_done_inst:in_conduit_0
	wire    [0:0] main_dpi_controller_inst_component_enabled_conduit;                                   // main_dpi_controller_inst:component_enabled -> split_component_start_inst:in_conduit
	wire          component_dpi_controller_streamer_inst_component_wait_for_stream_writes_conduit;      // component_dpi_controller_streamer_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_0
	wire          component_dpi_controller_streamer_inst_dpi_control_bind_conduit;                      // component_dpi_controller_streamer_inst:bind_interfaces -> streamer_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire          component_dpi_controller_streamer_inst_dpi_control_enable_conduit;                    // component_dpi_controller_streamer_inst:enable_interfaces -> streamer_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire          stream_sink_dpi_bfm_streamer_s_out_inst_dpi_control_stream_active_conduit;            // stream_sink_dpi_bfm_streamer_s_out_inst:stream_active -> streamer_component_dpi_controller_stream_active_concatenate_inst:in_conduit_0
	wire          concatenate_component_done_inst_out_conduit_conduit;                                  // concatenate_component_done_inst:out_conduit -> main_dpi_controller_inst:component_done
	wire          concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit;                // concatenate_component_wait_for_stream_writes_inst:out_conduit -> main_dpi_controller_inst:component_wait_for_stream_writes
	wire          streamer_component_dpi_controller_stream_active_concatenate_inst_out_conduit_conduit; // streamer_component_dpi_controller_stream_active_concatenate_inst:out_conduit -> component_dpi_controller_streamer_inst:stream_writes_active
	wire          split_component_start_inst_out_conduit_0_conduit;                                     // split_component_start_inst:out_conduit_0 -> component_dpi_controller_streamer_inst:component_enabled
	wire          streamer_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;     // streamer_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_streamer_s_in_inst:do_bind
	wire          streamer_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;   // streamer_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> stream_source_dpi_bfm_streamer_s_in_inst:enable
	wire          streamer_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;     // streamer_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> stream_sink_dpi_bfm_streamer_s_out_inst:do_bind
	wire          streamer_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;   // streamer_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> stream_sink_dpi_bfm_streamer_s_out_inst:enable
	wire          main_dpi_controller_inst_reset_ctrl_conduit;                                          // main_dpi_controller_inst:trigger_reset -> clock_reset_inst:trigger_reset
	wire          streamer_inst_return_valid;                                                           // streamer_inst:done -> component_dpi_controller_streamer_inst:done
	wire          component_dpi_controller_streamer_inst_component_return_stall;                        // component_dpi_controller_streamer_inst:stall -> streamer_inst:stall
	wire          clock_reset_inst_reset_reset;                                                         // clock_reset_inst:resetn -> [component_dpi_controller_streamer_inst:resetn, irq_mapper:reset, main_dpi_controller_inst:resetn, stream_sink_dpi_bfm_streamer_s_out_inst:resetn, stream_source_dpi_bfm_streamer_s_in_inst:resetn, streamer_inst:resetn]
	wire          component_dpi_controller_streamer_inst_component_irq_irq;                             // irq_mapper:sender_irq -> component_dpi_controller_streamer_inst:done_irq

	hls_sim_clock_reset #(
		.RESET_CYCLE_HOLD (4)
	) clock_reset_inst (
		.clock         (clock_reset_inst_clock_clk),                  //      clock.clk
		.resetn        (clock_reset_inst_reset_reset),                //      reset.reset_n
		.clock2x       (clock_reset_inst_clock2x_clk),                //    clock2x.clk
		.trigger_reset (main_dpi_controller_inst_reset_ctrl_conduit)  // reset_ctrl.conduit
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("streamer"),
		.COMPONENT_MANGLED_NAME       ("\\3fstreamer@@YAXXZ"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_AGENTS         (0),
		.COMPONENT_HAS_AGENT_RETURN   (0),
		.COMPONENT_NUM_OUTPUT_STREAMS (1)
	) component_dpi_controller_streamer_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                           //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                         //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                         //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_streamer_inst_dpi_control_bind_conduit),                      //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_streamer_inst_dpi_control_enable_conduit),                    //               dpi_control_enable.conduit
		.stream_writes_active             (streamer_component_dpi_controller_stream_active_concatenate_inst_out_conduit_conduit), // dpi_control_stream_writes_active.conduit
		.component_enabled                (split_component_start_inst_out_conduit_0_conduit),                                     //                component_enabled.conduit
		.component_done                   (component_dpi_controller_streamer_inst_component_done_conduit),                        //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_streamer_inst_component_wait_for_stream_writes_conduit),      // component_wait_for_stream_writes.conduit
		.agent_busy                       (),                                                                                     //                       agent_busy.conduit
		.read_implicit_streams            (),                                                                                     //            read_implicit_streams.conduit
		.readback_from_agents             (),                                                                                     //             readback_from_agents.conduit
		.start                            (component_dpi_controller_streamer_inst_component_call_valid),                          //                   component_call.valid
		.busy                             (streamer_inst_call_stall),                                                             //                                 .stall
		.done                             (streamer_inst_return_valid),                                                           //                 component_return.valid
		.stall                            (component_dpi_controller_streamer_inst_component_return_stall),                        //                                 .stall
		.done_irq                         (component_dpi_controller_streamer_inst_component_irq_irq),                             //                    component_irq.irq
		.returndata                       ()                                                                                      //                       returndata.data
	);

	tb_concatenate_component_done_inst concatenate_component_done_inst (
		.out_conduit  (concatenate_component_done_inst_out_conduit_conduit),           //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_streamer_inst_component_done_conduit)  // in_conduit_0.conduit
	);

	tb_concatenate_component_done_inst concatenate_component_wait_for_stream_writes_inst (
		.out_conduit  (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit),           //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_streamer_inst_component_wait_for_stream_writes_conduit)  // in_conduit_0.conduit
	);

	hls_sim_main_dpi_controller #(
		.NUM_COMPONENTS      (1),
		.COMPONENT_NAMES_STR ("streamer")
	) main_dpi_controller_inst (
		.clock                            (clock_reset_inst_clock_clk),                                            //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                          //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                          //                          clock2x.clk
		.component_enabled                (main_dpi_controller_inst_component_enabled_conduit),                    //                component_enabled.conduit
		.component_done                   (concatenate_component_done_inst_out_conduit_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit), // component_wait_for_stream_writes.conduit
		.trigger_reset                    (main_dpi_controller_inst_reset_ctrl_conduit)                            //                       reset_ctrl.conduit
	);

	tb_split_component_start_inst split_component_start_inst (
		.in_conduit    (main_dpi_controller_inst_component_enabled_conduit), //    in_conduit.conduit
		.out_conduit_0 (split_component_start_inst_out_conduit_0_conduit)    // out_conduit_0.conduit
	);

	hls_sim_stream_sink_dpi_bfm #(
		.COMPONENT_NAME                  ("streamer"),
		.INTERFACE_NAME                  ("@s_out"),
		.STREAM_DATAWIDTH                (352),
		.READY_LATENCY                   (0),
		.STREAM_BITSPERSYMBOL            (352),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_sink_dpi_bfm_streamer_s_out_inst (
		.clock              (clock_reset_inst_clock_clk),                                                         //                     clock.clk
		.resetn             (clock_reset_inst_reset_reset),                                                       //                     reset.reset_n
		.clock2x            (clock_reset_inst_clock2x_clk),                                                       //                   clock2x.clk
		.do_bind            (streamer_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),   //          dpi_control_bind.conduit
		.enable             (streamer_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit), //        dpi_control_enable.conduit
		.stream_active      (stream_sink_dpi_bfm_streamer_s_out_inst_dpi_control_stream_active_conduit),          // dpi_control_stream_active.conduit
		.sink_data          (streamer_inst_s_out_data),                                                           //                      sink.data
		.sink_ready         (streamer_inst_s_out_ready),                                                          //                          .ready
		.sink_valid         (streamer_inst_s_out_valid),                                                          //                          .valid
		.sink_startofpacket (1'b0),                                                                               //               (terminated)
		.sink_endofpacket   (1'b0),                                                                               //               (terminated)
		.sink_empty         (1'b0)                                                                                //               (terminated)
	);

	hls_sim_stream_source_dpi_bfm #(
		.COMPONENT_NAME                  ("streamer"),
		.INTERFACE_NAME                  ("@s_in"),
		.STREAM_DATAWIDTH                (352),
		.STREAM_BITSPERSYMBOL            (352),
		.EMPTY_WIDTH                     (0),
		.FIRST_SYMBOL_IN_HIGH_ORDER_BITS (0)
	) stream_source_dpi_bfm_streamer_s_in_inst (
		.clock        (clock_reset_inst_clock_clk),                                                         //              clock.clk
		.resetn       (clock_reset_inst_reset_reset),                                                       //              reset.reset_n
		.clock2x      (clock_reset_inst_clock2x_clk),                                                       //            clock2x.clk
		.do_bind      (streamer_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),   //   dpi_control_bind.conduit
		.enable       (streamer_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // dpi_control_enable.conduit
		.source_data  (stream_source_dpi_bfm_streamer_s_in_inst_source_data),                               //             source.data
		.source_ready (stream_source_dpi_bfm_streamer_s_in_inst_source_ready),                              //                   .ready
		.source_valid (stream_source_dpi_bfm_streamer_s_in_inst_source_valid)                               //                   .valid
	);

	tb_streamer_component_dpi_controller_bind_conduit_fanout_inst streamer_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_streamer_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (streamer_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (streamer_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_streamer_component_dpi_controller_bind_conduit_fanout_inst streamer_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_streamer_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (streamer_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (streamer_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_concatenate_component_done_inst streamer_component_dpi_controller_stream_active_concatenate_inst (
		.out_conduit  (streamer_component_dpi_controller_stream_active_concatenate_inst_out_conduit_conduit), //  out_conduit.conduit
		.in_conduit_0 (stream_sink_dpi_bfm_streamer_s_out_inst_dpi_control_stream_active_conduit)             // in_conduit_0.conduit
	);

	tb_streamer_inst streamer_inst (
		.start       (component_dpi_controller_streamer_inst_component_call_valid),   //   call.valid
		.busy        (streamer_inst_call_stall),                                      //       .stall
		.clock       (clock_reset_inst_clock_clk),                                    //  clock.clk
		.resetn      (clock_reset_inst_reset_reset),                                  //  reset.reset_n
		.done        (streamer_inst_return_valid),                                    // return.valid
		.stall       (component_dpi_controller_streamer_inst_component_return_stall), //       .stall
		.s_in_data   (stream_source_dpi_bfm_streamer_s_in_inst_source_data),          //   s_in.data
		.s_in_ready  (stream_source_dpi_bfm_streamer_s_in_inst_source_ready),         //       .ready
		.s_in_valid  (stream_source_dpi_bfm_streamer_s_in_inst_source_valid),         //       .valid
		.s_out_data  (streamer_inst_s_out_data),                                      //  s_out.data
		.s_out_ready (streamer_inst_s_out_ready),                                     //       .ready
		.s_out_valid (streamer_inst_s_out_valid)                                      //       .valid
	);

	tb_irq_mapper irq_mapper (
		.clk        (clock_reset_inst_clock_clk),                               //       clk.clk
		.reset      (~clock_reset_inst_reset_reset),                            // clk_reset.reset
		.sender_irq (component_dpi_controller_streamer_inst_component_irq_irq)  //    sender.irq
	);

endmodule
