// soc_system_streamer_0.v

// Generated using ACDS version 21.1 850

`timescale 1 ps / 1 ps
module soc_system_streamer_0 (
		input  wire         avs_tuple_in_read,        //  avs_tuple_in.read
		output wire [511:0] avs_tuple_in_readdata,    //              .readdata
		input  wire         avs_tuple_in_write,       //              .write
		input  wire [511:0] avs_tuple_in_writedata,   //              .writedata
		input  wire         avs_tuple_in_address,     //              .address
		input  wire [63:0]  avs_tuple_in_byteenable,  //              .byteenable
		input  wire         avs_tuple_out_read,       // avs_tuple_out.read
		output wire [511:0] avs_tuple_out_readdata,   //              .readdata
		input  wire         avs_tuple_out_write,      //              .write
		input  wire [511:0] avs_tuple_out_writedata,  //              .writedata
		input  wire         avs_tuple_out_address,    //              .address
		input  wire [63:0]  avs_tuple_out_byteenable, //              .byteenable
		input  wire         clock,                    //         clock.clk
		input  wire         resetn                    //         reset.reset_n
	);

	streamer_internal streamer_internal_inst (
		.clock                    (clock),                    //         clock.clk
		.resetn                   (resetn),                   //         reset.reset_n
		.avs_tuple_in_read        (avs_tuple_in_read),        //  avs_tuple_in.read
		.avs_tuple_in_readdata    (avs_tuple_in_readdata),    //              .readdata
		.avs_tuple_in_write       (avs_tuple_in_write),       //              .write
		.avs_tuple_in_writedata   (avs_tuple_in_writedata),   //              .writedata
		.avs_tuple_in_address     (avs_tuple_in_address),     //              .address
		.avs_tuple_in_byteenable  (avs_tuple_in_byteenable),  //              .byteenable
		.avs_tuple_out_read       (avs_tuple_out_read),       // avs_tuple_out.read
		.avs_tuple_out_readdata   (avs_tuple_out_readdata),   //              .readdata
		.avs_tuple_out_write      (avs_tuple_out_write),      //              .write
		.avs_tuple_out_writedata  (avs_tuple_out_writedata),  //              .writedata
		.avs_tuple_out_address    (avs_tuple_out_address),    //              .address
		.avs_tuple_out_byteenable (avs_tuple_out_byteenable)  //              .byteenable
	);

endmodule
