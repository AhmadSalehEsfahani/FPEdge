// soc_system_streamer_0.v

// Generated using ACDS version 21.1 850

`timescale 1 ps / 1 ps
module soc_system_streamer_0 (
		input  wire        avs_cra_read,       // avs_cra.read
		output wire [63:0] avs_cra_readdata,   //        .readdata
		input  wire        avs_cra_write,      //        .write
		input  wire [63:0] avs_cra_writedata,  //        .writedata
		input  wire [3:0]  avs_cra_address,    //        .address
		input  wire [7:0]  avs_cra_byteenable, //        .byteenable
		input  wire        clock,              //   clock.clk
		output wire        done_irq,           //     irq.irq
		input  wire        resetn              //   reset.reset_n
	);

	streamer_internal streamer_internal_inst (
		.clock              (clock),              //   clock.clk
		.resetn             (resetn),             //   reset.reset_n
		.done_irq           (done_irq),           //     irq.irq
		.avs_cra_read       (avs_cra_read),       // avs_cra.read
		.avs_cra_readdata   (avs_cra_readdata),   //        .readdata
		.avs_cra_write      (avs_cra_write),      //        .write
		.avs_cra_writedata  (avs_cra_writedata),  //        .writedata
		.avs_cra_address    (avs_cra_address),    //        .address
		.avs_cra_byteenable (avs_cra_byteenable)  //        .byteenable
	);

endmodule
