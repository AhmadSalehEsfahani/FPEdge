// tb_streamer_inst.v

// Generated using ACDS version 21.1 850

`timescale 1 ps / 1 ps
module tb_streamer_inst (
		input  wire         start,       //   call.valid
		output wire         busy,        //       .stall
		input  wire         clock,       //  clock.clk
		input  wire         resetn,      //  reset.reset_n
		output wire         done,        // return.valid
		input  wire         stall,       //       .stall
		input  wire [351:0] s_in_data,   //   s_in.data
		output wire         s_in_ready,  //       .ready
		input  wire         s_in_valid,  //       .valid
		output wire [351:0] s_out_data,  //  s_out.data
		input  wire         s_out_ready, //       .ready
		output wire         s_out_valid  //       .valid
	);

	streamer_internal streamer_internal_inst (
		.clock       (clock),       //  clock.clk
		.resetn      (resetn),      //  reset.reset_n
		.s_in_data   (s_in_data),   //   s_in.data
		.s_in_ready  (s_in_ready),  //       .ready
		.s_in_valid  (s_in_valid),  //       .valid
		.s_out_data  (s_out_data),  //  s_out.data
		.s_out_ready (s_out_ready), //       .ready
		.s_out_valid (s_out_valid), //       .valid
		.start       (start),       //   call.valid
		.busy        (busy),        //       .stall
		.done        (done),        // return.valid
		.stall       (stall)        //       .stall
	);

endmodule
